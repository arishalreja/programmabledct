library IEEE;
use IEEE.STD_LOGIC_1164.all;

package mem_content is

-- content of m_0_0
constant m_0_0_0 : BIT_VECTOR := X"C49324C144C0F3F32B0994ABB1A49946D92AFBD2E499000500010000080006D8";
constant m_0_0_1 : BIT_VECTOR := X"3D484000008C79DAAACA49A248BDE4C550FED992CE14CE1F3B9F995856C9B8AF";
constant m_0_0_2 : BIT_VECTOR := X"BEEF2673DF4C6455448448449401128600DD5E0C976930800001FA68EF0E0FFB";
constant m_0_0_3 : BIT_VECTOR := X"1C79C5674A32F2B39DE71971BB18749249328951692A5D091612124A3AD45547";
constant m_0_0_4 : BIT_VECTOR := X"7CB23FDFFD5BFFD5AA5FFEAD447FFAB5019BBED52FFDD5F2099A8D485B6BB6A3";
constant m_0_0_5 : BIT_VECTOR := X"1A999AADED9BDB7E3C2C87F7FECF6FFECF7BDB97FF67BDED8BFFB3DEF9747FF7";
constant m_0_0_6 : BIT_VECTOR := X"6854972B5277C7A4003C3ADD6D2DCD15F18B5DD5E15659B6EFA4B6B57BEBDD5E";
constant m_0_0_7 : BIT_VECTOR := X"F3FF26EA48480669FB7EDFB7EDFB5FD7F77B5EF6F7ED5497209DF9E000F0DABF";
constant m_0_0_8 : BIT_VECTOR := X"771212F3FF06EA484904BCFFC1BAB21212F09BD49BA12F3FF06EAC84943E9212";
constant m_0_0_9 : BIT_VECTOR := X"ECA2BBD94537B28AEF6514DECA2BBD94537B28AEF652E2B7B38A55EB674AA742";
constant m_0_0_A : BIT_VECTOR := X"95A7F5E0A5487F683754BF25583FED26EA9521B5FED80277C5A8A128AEF6514D";
constant m_0_0_B : BIT_VECTOR := X"D77D266D55B8B316F0DFD81DA5FFF81FFFCE7F67AFDDD9999762ED8EC59B15DB";
constant m_0_0_C : BIT_VECTOR := X"4EFDFA99F39BE6607021F9DF9EA6EDCAC249598B2C960C6FFFFBDFA3E597BF7A";
constant m_0_0_D : BIT_VECTOR := X"0000000000000000000000000000000001E243A027FBE2E7DF37532E66F3BF3E";
constant m_0_0_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000002000";

-- content of m_0_1
constant m_0_1_0 : BIT_VECTOR := X"488E3389239716B6268F601CBF78F40B9B1051846273020203020000080005B8";
constant m_0_1_1 : BIT_VECTOR := X"0DC550000092D67EF9A0541876046400CF5ADB233892397168B7B1346D0F641C";
constant m_0_1_2 : BIT_VECTOR := X"8E23A3104646A20E3B66A67B555BA89C00DBF5551AAA5C5000016997BAA28916";
constant m_0_1_3 : BIT_VECTOR := X"248B66D9DA50D36CB6E905D851869FB1089AD12C29810FCCC391196B52438EB0";
constant m_0_1_4 : BIT_VECTOR := X"548A93452D3052D320429699010A5A64449CAD232525737E0F773FC57E23801D";
constant m_0_1_5 : BIT_VECTOR := X"2F0A8C6203045C2290E304D14A6AA14A6AB2A8B0A535594448529AACA9050A52";
constant m_0_1_6 : BIT_VECTOR := X"05A133203CD570F00001DD2E97A09260320FEC7AD2F13A802BD1890E0AF3C7AD";
constant m_0_1_7 : BIT_VECTOR := X"ADEFCDA627267ABF5A73B5A73B5A7395AF3B4A72F7D208116A15787400077F76";
constant m_0_1_8 : BIT_VECTOR := X"55EDC2ADEFCDA6272770AB7BFB688DEDC2AE4DD3369C2ADEFCDA237B13C88DC2";
constant m_0_1_9 : BIT_VECTOR := X"1653722CA6E4594D48B29A91653722CA6E4594D48B2A336458A52AD511BFDDF8";
constant m_0_1_A : BIT_VECTOR := X"1FBAD75481C52D4B245037455565A9648A0714B4BD2B7855FA54DED4D48B29A9";
constant m_0_1_B : BIT_VECTOR := X"F28122ED401E341EB2024BB7A4206BB7E5CBA869CFC578C983E7E7A7CF8F478F";
constant m_0_1_C : BIT_VECTOR := X"1D4ED413A9D512A052C403ED682F56E7500A08E3041F95200003A96A514753F0";
constant m_0_1_D : BIT_VECTOR := X"00000000000000000000000000000000015E2AADBC7DAA53A95282657D47DBB5";
constant m_0_1_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_2
constant m_0_2_0 : BIT_VECTOR := X"C6688A047A1C489888A44650D80205701488B8C8B6440000000100000FFFFA58";
constant m_0_2_1 : BIT_VECTOR := X"44245000008B1C488229347516927612AC485C18A147A0C48A44C44511A44650";
constant m_0_2_2 : BIT_VECTOR := X"6E9BB99D377338E991351340040D01F000CD4700C00882400001200283806008";
constant m_0_2_3 : BIT_VECTOR := X"146451110025288A45E2C72476C6F94FA68DE44D97A340A2D94D45178426287A";
constant m_0_2_4 : BIT_VECTOR := X"245E58508C3508C355284618B8A1186AE2E87C89C883C930E008440C4816CD69";
constant m_0_2_5 : BIT_VECTOR := X"48A2009750F2A685C3967E1422E41422E419054A11720C92B508B90640A8A117";
constant m_0_2_6 : BIT_VECTOR := X"44D4B322224F3C45FFFF388C46C808C451FD82E85C0B32041E645D42C79C2E85";
constant m_0_2_7 : BIT_VECTOR := X"5BB489A57ED42442102108484200A4014802048161DADCB36493EF4BFFFCEC66";
constant m_0_2_8 : BIT_VECTOR := X"4F90935BB489A57ED524D6ED2A697B90935DA952A68935BB4A9A5EE44B9CC893";
constant m_0_2_9 : BIT_VECTOR := X"8309790612F20C25E4184BC8309590612B20C256418609720CF0F1830E190C92";
constant m_0_2_A : BIT_VECTOR := X"C3AE4070880C6401801113319C4C8010022031D8DDA8924F93425902564184AC";
constant m_0_2_B : BIT_VECTOR := X"4103A8668B5192F10A8845845584418480C872103903C717871E104E1C609428";
constant m_0_2_C : BIT_VECTOR := X"300008AE00A8AABFC88806448440204001AAEA01B7F82040000644A528888955";
constant m_0_2_D : BIT_VECTOR := X"00000000000000000000000000000000012063D90288840C000115C0A22C8800";
constant m_0_2_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000006000";

-- content of m_0_3
constant m_0_3_0 : BIT_VECTOR := X"A10B42C202C023834395C40131B11D40C1880000045C01010101000000000289";
constant m_0_3_1 : BIT_VECTOR := X"9C01D000004044923CF0842084087000081215842C202D02B91C1A1C8715C401";
constant m_0_3_2 : BIT_VECTOR := X"4F4381008702004019A19A1996CA66F600081164022C10180000499A28B60334";
constant m_0_3_3 : BIT_VECTOR := X"8A11C8726D0804391CF085085486E51A10880208100200908021212008040051";
constant m_0_3_4 : BIT_VECTOR := X"490804488BB088BB000445DA001117680000A8804885442201140C4593000428";
constant m_0_3_5 : BIT_VECTOR := X"08C465A2204603120BA379122209C22209C270A11104E1280088827096121110";
constant m_0_3_6 : BIT_VECTOR := X"42D4956217959325FFFF2080410808055576C54C081104042B0488000A8854C0";
constant m_0_3_7 : BIT_VECTOR := X"AFB699AAACD4E89EE71CC731CC63B9E7718CE31CAC9ADC9529E54493FFFCB70C";
constant m_0_3_8 : BIT_VECTOR := X"9535BDAFB6B9AAACD4EF6BEDA66AAB35BDA8895666BBDAFB699AAACD2B4F85BD";
constant m_0_3_9 : BIT_VECTOR := X"394542728A84E51509CA2A1394542728A84E51509CA2C544E594F8F164884437";
constant m_0_3_A : BIT_VECTOR := X"13F89116D345C91A0CDA67E155C923619B4D176E09A1379533515351589CA2B1";
constant m_0_3_B : BIT_VECTOR := X"24A30CF5010C92E766845959D1445D5924EB2201B2454869C43244C864C99099";
constant m_0_3_C : BIT_VECTOR := X"F3366C4CDECCE0DFBCCC0466C64B3168A1C3832D2BE73108000622E5B25844C9";
constant m_0_3_D : BIT_VECTOR := X"0000000000000000000000000000000000722D718B8CCCB46645898B333CCDDB";
constant m_0_3_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000004000";

-- content of m_0_4
constant m_0_4_0 : BIT_VECTOR := X"28040110C10004241C020421025020511608A010842207020302000007FFF811";
constant m_0_4_1 : BIT_VECTOR := X"C010800000521080110000A00180380000005220100C1100402120E038020021";
constant m_0_4_2 : BIT_VECTOR := X"0701C120038241531925925916C9640800010424220185080000008002125100";
constant m_0_4_3 : BIT_VECTOR := X"AA820382204A01C020F0110110B00162000A00C30462C4803000002802040040";
constant m_0_4_4 : BIT_VECTOR := X"1B01000282082820A2814105100504145000228408C104021100C00081001400";
constant m_0_4_5 : BIT_VECTOR := X"9CC440810652531088000000A1E340A1E358D00050F1AC68002878D63210050F";
constant m_0_4_6 : BIT_VECTOR := X"426DB76A17849324000000C0400C0805550000244180941409040499424A0244";
constant m_0_4_7 : BIT_VECTOR := X"0092541881D3A508D631AD631AD610A4214AC6B08DBA65B765E124C80000250D";
constant m_0_4_8 : BIT_VECTOR := X"84743C0092741881D28F0024950600743C0283055023C0092541801D095A843C";
constant m_0_4_9 : BIT_VECTOR := X"682018D04031A080634100C682018D04031A08063417A031A00245AB465B2D87";
constant m_0_4_A : BIT_VECTOR := X"31C000029800800844130381108001088260024A1BA4878483C807480634100C";
constant m_0_4_B : BIT_VECTOR := X"F3A02AB0A114820054C014201014342000E8830800010405C712244E04489C58";
constant m_0_4_C : BIT_VECTOR := X"57EEDC39BBDD82A000CC02FDCC3FF4EA104A4AA42C0035600002FDC77BD1FBB5";
constant m_0_4_D : BIT_VECTOR := X"0000000000000000000000000000000000000E01AE1FBB70FDDB87377765FBB7";
constant m_0_4_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000002000";

-- content of m_0_5
constant m_0_5_0 : BIT_VECTOR := X"A050141054128808080414A3240441140422AA52908401010000000007FFF815";
constant m_0_5_1 : BIT_VECTOR := X"5149900000405192320A28AA28A2B2851292C4014105402880404040104414A3";
constant m_0_5_2 : BIT_VECTOR := X"5715950A2B2A145155215215068854E00009142091098488000049522A340AA0";
constant m_0_5_3 : BIT_VECTOR := X"8A040106680290804070040A44046540452AA85145285085140A0A2AA2915114";
constant m_0_5_4 : BIT_VECTOR := X"1D22A08250422504085128205144A08105228254025410200880C15092483282";
constant m_0_5_5 : BIT_VECTOR := X"0A111220A1080848A720F82095E34895E358D2144AF1AC795A2578D6365344AF";
constant m_0_5_6 : BIT_VECTOR := X"BA100C09505044A1FFFEA251290545111472541128545532A080A28528214112";
constant m_0_5_7 : BIT_VECTOR := X"A249325A8928A458D6B1AC6358D6B58C635AC6318425100C00141523FFFA9281";
constant m_0_5_8 : BIT_VECTOR := X"504A02A249325A892980A8924C96A24A02A3708CC9602A249325A89285261202";
constant m_0_5_9 : BIT_VECTOR := X"6880B8D10171A202E34405C6880B8D10171A202E344180B1A2081060D5008040";
constant m_0_5_A : BIT_VECTOR := X"25C095060A51C9502A8147A451992A05502947254250005044A024A02E34405C";
constant m_0_5_B : BIT_VECTOR := X"4920017414B010E54C50B441151290412AC28942B25410A19154A946A1028D12";
constant m_0_5_C : BIT_VECTOR := X"42A54A08928A903F94000054A512AA49044040551FE50250000054B52290A951";
constant m_0_5_D : BIT_VECTOR := X"0000000000000000000000000000000000528F20124A952254A9411222A0A952";
constant m_0_5_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_6
constant m_0_6_0 : BIT_VECTOR := X"2A91A4556454D111A968945B1896890650AA9392A68900000000000007FFF859";
constant m_0_6_1 : BIT_VECTOR := X"D90480000052118104534A134AB4B4A6D480D8AA4556454D16888D4B5268945B";
constant m_0_6_2 : BIT_VECTOR := X"97A5A5134B4A252D5981981996E066020025046E8664B458000005980217033A";
constant m_0_6_3 : BIT_VECTOR := X"AAA8B5262248DA968AF0A1401401000B6928CD5551AB54A95552D28328D66D66";
constant m_0_6_4 : BIT_VECTOR := X"19A02AB4964349642A1A4B2140692C85012A049442901497433A59018168A482";
constant m_0_6_5 : BIT_VECTOR := X"02DDDA80A14B4B6A340082AD24E36D24E378DA069271BC7D534938DE37426927";
constant m_0_6_6 : BIT_VECTOR := X"4A56D5B2534050A6000022914809A9D775801115A84441A480A622042021115A";
constant m_0_6_7 : BIT_VECTOR := X"024932488A498108529484214A4210842158C6B1AEC956D5B4D01028000080A6";
constant m_0_6_8 : BIT_VECTOR := X"40929A024932488A49A680924C9222929A0490A4C929A024932488A4D4AA0A9A";
constant m_0_6_9 : BIT_VECTOR := X"6EAA98DD5531BAAA637554C6EAA98DD5531BAAA63752AAB1BAAA54A94148A453";
constant m_0_6_A : BIT_VECTOR := X"05C80442DB00805D0CDB638510900B819B6C02010C949340512AA92AA637554C";
constant m_0_6_B : BIT_VECTOR := X"6DE105F28534CB00049A908805A4B0880AC88A6A801014A59744890A89121502";
constant m_0_6_C : BIT_VECTOR := X"53366DAEDAECD06004660066D65B337DD9014164BC011BD8000066E5B2F0CDD9";
constant m_0_6_D : BIT_VECTOR := X"0000000000000000000000000000000000100608DB0CD9B866CDB5DBBB34CD9B";
constant m_0_6_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000002000";

-- content of m_0_7
constant m_0_7_0 : BIT_VECTOR := X"0042109050920A0A0A4504200520504081000840101101010101000000000241";
constant m_0_7_1 : BIT_VECTOR := X"D00080000002000102882288208232210200050108050820A450505214050020";
constant m_0_7_2 : BIT_VECTOR := X"47119008232011110420420426281004002400220100800800000550001502A0";
constant m_0_7_3 : BIT_VECTOR := X"00052140000800A4527480080480011004002041002040041008888080011010";
constant m_0_7_4 : BIT_VECTOR := X"0100002240002400020120001004800040000240004000910080401080001200";
constant m_0_7_5 : BIT_VECTOR := X"0000000020414002000000089080409080401080484020080024201006020484";
constant m_0_7_6 : BIT_VECTOR := X"2202449910001022000080402044440114800000000000120002000000000000";
constant m_0_7_7 : BIT_VECTOR := X"20003008012181085294A52908421084214A5210A42402449000000000020021";
constant m_0_7_8 : BIT_VECTOR := X"0048002000300801218008000C02204800224024C02002000300881200020000";
constant m_0_7_9 : BIT_VECTOR := X"0800201000402000804001008002010004020008040080002000002040000000";
constant m_0_7_A : BIT_VECTOR := X"01C800421A1080150A8343A0108002A150684200024000000480048008040010";
constant m_0_7_B : BIT_VECTOR := X"4920017280844901044014504012145000C08000000000018100000200000400";
constant m_0_7_C : BIT_VECTOR := X"52A54A0892AA800000220254A412AA490040004488010A50000054852290A911";
constant m_0_7_D : BIT_VECTOR := X"0000000000000000000000000000000000008408520A952854A94112AAA4A952";
constant m_0_7_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_0
constant m_1_0_0 : BIT_VECTOR := X"0000000000000000000000080000000000000000000000000000000000000000";
constant m_1_0_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_2 : BIT_VECTOR := X"302B550056AA53E19B235C46394F880140807C6803C2802A2C00000000000000";
constant m_1_0_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000724AC77CE";
constant m_1_0_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_1
constant m_1_1_0 : BIT_VECTOR := X"0000000000000000000000080000000000000000000000000000000000000000";
constant m_1_1_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_2 : BIT_VECTOR := X"104C660098CC30608537586EB0C1B8017180675801F380675800000000000000";
constant m_1_1_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000601988A0C";
constant m_1_1_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_2
constant m_1_2_0 : BIT_VECTOR := X"0000000000000000000000180000000000000000000000000000000000000000";
constant m_1_2_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_2 : BIT_VECTOR := X"58707800E0F051ABA26E02DC054688011000704803B280092C00000000000000";
constant m_1_2_3 : BIT_VECTOR := X"00000000000000000000000000000000000000000000000000000000B8DDF4C1";
constant m_1_2_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_3
constant m_1_3_0 : BIT_VECTOR := X"0000000000000000000000180000000000000000000000000000000000000000";
constant m_1_3_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_2 : BIT_VECTOR := X"1A01800403001930A86610CC2064C00120007868019200230600000000000000";
constant m_1_3_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000414BCA048";
constant m_1_3_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_4
constant m_1_4_0 : BIT_VECTOR := X"0000000000000000000000080000000000000000000000000000000000000000";
constant m_1_4_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_2 : BIT_VECTOR := X"0301FF8603FF247B05184A309491F80161000F10045780777800000000000000";
constant m_1_4_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000281410E05";
constant m_1_4_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_5
constant m_1_5_0 : BIT_VECTOR := X"0000000000000000000000080000000000000000000000000000000000000000";
constant m_1_5_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_2 : BIT_VECTOR := X"F37FFF8203FF7FDBFF7FFEFFFDFF6804008009000200802A2A00000000000000";
constant m_1_5_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000779F9FF9E";
constant m_1_5_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_6
constant m_1_6_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_2 : BIT_VECTOR := X"7A7E0004FC007FFBBF7F1EFE3DFFE80010800808000080020A00000000000000";
constant m_1_6_3 : BIT_VECTOR := X"00000000000000000000000000000000000000000000000000000007BDFDFFCF";
constant m_1_6_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_7
constant m_1_7_0 : BIT_VECTOR := X"0000000000000000000000080000000000000000000000000000000000000000";
constant m_1_7_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_2 : BIT_VECTOR := X"00000000000000000000000000000000800000000202000A0000000000000000";
constant m_1_7_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";


end mem_content;

package body mem_content is

end mem_content;

