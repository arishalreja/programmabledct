-- This module is a wrapper that creates the Wishbone logic around the DCT core
-- and the Output buffer

library ieee;
use ieee.std_logic_1164.all;

library WORK;
use WORK.MDCT_PKG.all;
use IEEE.NUMERIC_STD.all;
use WORK.dpmem;

 entity WBOPRT08 is
   port(
-- WISHBONE SLAVE interface for DCT acc core:
   ACK_O: out std_logic;  -- WBC Acknowledge Output signal
   CLK_I: in std_logic;   -- WBC Clock signal
   DAT_I: in std_logic_vector( 7 downto 0 ); -- 8 bit WBC Data input bus
   DAT_O: out std_logic_vector( 7 downto 0 );-- 8 bit WBC Data output bus
   RST_I: in std_logic; -- WBC Reset In signal
   STB_I: in std_logic; -- WBC Strobe In signal
   CYC_I : in std_logic; -- WBC Cycle In signal
   WE_I: in std_logic -- WBC Write Enable In signal
   );
 end entity WBOPRT08;

 architecture WBOPRT081 of WBOPRT08 is

component MDCT_comp IS	 -- This component is the original non WBC DCT core
	port   (	  
		clk          : in STD_LOGIC;  
		rst          : in std_logic;
      dcti         : in std_logic_vector(IP_W-1 downto 0);
      idv          : in STD_LOGIC;

      odv          : out STD_LOGIC;
      dcto         : out std_logic_vector(COE_W-1 downto 0);
      odv1         : out STD_LOGIC;
      dcto1        : out std_logic_vector(OP_W-1 downto 0)
      );
      end component MDCT_comp; 
  
  FOR ALL:  MDCT_comp USE ENTITY WORK.MDCT(RTL);
    
 component dpmem_comp IS -- This component is the Output Buffer
   port  (
      clk          : in STD_LOGIC;
      reset        : in STD_LOGIC;
      empty	   : out STD_LOGIC; -- cclin
      Data_In  : in  std_logic_vector(15 DOWNTO 0);    -- input data
      Data_Out : out std_logic_vector(7 DOWNTO 0);    -- output Data
      WR          : in  std_logic;                                -- Write Enable
      RE          : in  std_logic                                 -- Read Enable
      );
  end component dpmem_comp;
  
   FOR ALL: dpmem_comp USE ENTITY WORK.dpmem(dpmem_v1);                               
    
   signal Q: std_logic_vector( 15 downto 0 ); -- The 16 bit extended version of the 12 
                                              -- bit DCT core output
   signal R: std_logic_vector( 7 downto 0); -- This signal is mapped to the 8 bit output
                                            -- of the wrapper, output of the Output Buffer
   signal S: std_logic_vector( 15 downto 0); -- This forms the input to the output buffer
   signal odvtemp: STD_LOGIC;
   signal idvtemp: STD_LOGIC;
   signal odv1temp: STD_LOGIC;
   signal Data_Intemp: std_logic_vector(7 downto 0);
   signal WRtemp: STD_LOGIC;
   signal REtemp: STD_LOGIC;
   signal dcto1temp: std_logic_vector(OP_W-1 downto 0);
   signal flag1: STD_LOGIC;  -- This is used to ensure that no data is read
                             -- from the mem buf until it contains the first
                             -- new output data value data
--   signal  All_Outs     : out std_logic;
   --cclin
   signal empty: STD_LOGIC;
   signal ack_tmp: STD_LOGIC;
    
   begin
      REG: process( CLK_I )
    VARIABLE count : INTEGER := 0; 
         begin
           -- The following logic handles the control logic for the WBC interface            
           if ( falling_edge( CLK_I ) ) then 

	-- masked by cclin
              --if ((odvtemp and flag1) = '1') then  -- If there is output data to be read
              --    REtemp <= '1'; -- Read enable (for the buffer) is set
              --end if;  
              
              if (odvtemp = '1') then -- If data is being written to output buffer
                                      -- during the next rising edge
                  flag1 <= '1';  -- Set flag
              else
                  flag1 <= '0';  -- else null it          
              end if;
              
              if (REtemp = '1') then    -- if read is enabled, the next rising edge
                                        -- there will be data in R
                  count := count + 1;   -- Increment counter
                  --ACK_O <= ((STB_I and (not(WE_I)))); -- Ack = STB.(WE)'
              else                          
                  --ACK_O <= ((STB_I) and (WE_I));   -- Ack = STB.WE    
              end if;
              
              if (count = 129) then       -- End of read (no more read)      
                  count := 0;             -- Reset Counter
              --    REtemp <= '0';          -- Read Enable nulled
              end if;
              -- Note - Reset operation is taken care of internally.
              --DAT_O <= R; -- The output of the Output buffer is written to DAT_O via R every falling edge     
              S <= Q; -- The sign extended output of the DCT core
                      -- is written to the Output buffer            
            end if; 
             
      end process REG;
   
   idvtemp <= STB_I and WE_I;

   --cclin
   DAT_O <= R; 
   REtemp	<= (not empty) and STB_I and (not WE_I);
   ACK_O	<= ack_tmp;
   process ( REtemp, WE_I, STB_I, ack_tmp) begin
      if (REtemp = '1') then    
          ack_tmp <= ((STB_I and (not(WE_I)))); -- Ack = STB.(WE)'
      else                          
          ack_tmp <= ((STB_I) and (WE_I));   -- Ack = STB.WE    
      end if;
   end process;
   
   Q(15) <= Q(11); -- The 12 bit output of the DCT is extended to 16 bits
   Q(14) <= Q(11); -- by logical sign extension
   Q(13) <= Q(11);
   Q(12) <= Q(11);
   
   YOT1: MDCT_comp 
   PORT MAP(
   clk => CLK_I,
   rst => RST_I,
   dcti => DAT_I,
   idv => idvtemp,
   odv => odvtemp,
   dcto => Q (11 downto 0),-- The DCT core writes its 12 bit output to the Q signal
   odv1 => odv1temp,
   dcto1 => dcto1temp);
   
   YOT2: dpmem_comp
   PORT MAP(
   clk		=> CLK_I,
   reset	=> RST_I,
   empty	=> empty, --cclin
   Data_In	=> S,  -- The S signal feeds the input to the output buffer
   Data_Out	=> R, -- The Output buffer writes its data to the R signal
   WR		=> odvtemp,
   RE		=> REtemp);
  -- All_Out => All_Outs);

end architecture WBOPRT081;
  
   

